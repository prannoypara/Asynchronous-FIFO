`timescale 1ns / 1ps

module tb_async_fifo;
reg wr_clk,rd_clk,reset;
wire wr_full,rd_empty;
wire [7:0] data_out;

async_fifo uut(data_out, wr_full, rd_empty,rd_clk, wr_clk, reset);


initial 
begin
wr_clk=0;
rd_clk=0;
reset=1;

end


initial
#5 reset=0;

always
#50 wr_clk=~wr_clk; //freq=10MHz

always
#500 rd_clk=~rd_clk; //freq= 1MHz

endmodule
